� �  �                      * * * * * * * * * * * * * * * * * * *                                           * p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p*                                           * p p p p pSpUpPpEpRpBpIpLpLp'pSp pRpEpSpTpApUpRpApNpTp p p p p p p p p*                                           * p p p p p p p p p pBprpepapkpfpapsptp pMpepnpup p p p p p p p p p p p*                                           * p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p*                                           * p p p p p p1p)pCprpepapmpepdp pSpiplpipcpopnp pCphpipppsp.p.p.p p p p*                                           * p p p p p p p pSptpoppp pBpepfpoprpep pIpcpep pCprpepapmp!p p p p p p*                                           * p p p p p p2p)pFprpipepdp pCpiprpcpupiptpsp.p.p.p p p p p p p p p p p*                                           * p p p p p p p pTpipmpep pTpop pWpapkpep-pUppp!p p p p p p p p p p p p*                                           * p p p p p p3p)pSpcprpapmpbplpepdp pDpipspkpeptptpepsp p p p p p p p p*                                           * p p p p p p p pSpupnpnpyp-pSpipdpep pUppp!p p p p p p p p p p p p p p*                                           * p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p*                                           * * * * * * * * * * * * * * * * * * *                                                                                                                                                                                                                                                                              It's similar to choosing breakfast at your favorite restaurant.             <!> Please place your order by pressing the number key                              corresponding to your choice:                                                                                                                                   Or Press Escape To Exit This Demo...                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   � �  �