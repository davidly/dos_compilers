� �  �     ` `  ` `     ` ` ` !p p @p p #p p $p p %p p ^p p &p p *p p (p p )p p _p p +p p  ` ` ` ` ` ` ` `  `N`u`m` ` S`c`r`o`l`l`          F`1` F`2`    E`s`c` 1p p 2p p 3p p 4p p 5p p 6p p 7p p 8p p 9p p 0p p -p p =p p  ` ``�`�` ` ` `  `L`o`c`k`  `L`o`c`k` `                                                                           `B`r`e`a`k`           ` `  ` `    �``�` ` ` Qp p Wp p Ep p Rp p Tp p Yp p Up p Ip p Op p Pp p {p p  p}p p  ` ` ` ` ` 7p p 8p p 9p p �a�a�a          F`3` F`4`     `�``�` `  p p  p p  p p  p p  p p  p p  p p  p p  p p  p p [p p  p]p p  ` ` ` ` `  p p p p  p p -` ` `                                                               ` `�` ` `                        ` `  ` `     ` ` ` ` ` ` Ap p Sp p Dp p Fp p Gp p Hp p Jp p Kp p Lp p :p p "p p ~p p  ``�` ` ` 4p p 5p p 6p p  f f `          F`5` F`6`     `C`t`r`l` `  p p  p p  p p  p p  p p  p p  p p  p p  p p ;p p 'p p `p p  ` ` ` ` ` p�p  p p �pp  ` ` `                                                                              ` ` `           ` `  ` `     `/`\` ` |p p Zp p Xp p Cp p Vp p Bp p Np p Mp p <p p >p p ?p p  `/`\` ` P`r`t`S`c` 1p p 2p p 3p p  ` ` `          F`7` F`8`     `�`�` ` \p p  p p  p p  p p  p p  p p  p p  p p ,p p .p p /p p  `�`�` ` *` ` ` ` `  p p p p  p p +` ` `                                                                              ` ` `           ` `  ` ` `    ` ` ` ` ` ` ` ۗۗۗۗۗۗۗۗۗۗۗۗۗۗۗۗۗۗۗۗۗۗۗۗۗۗۗۗ  ` `C`a`p`s` ` `  p0p p p w  w.p p p w  ` ` `          F`9` F`1`0`    ` `A`l`t` ` ` ۗۗۗۗۗۗۗۗۗۗۗۗۗۗۗۗۗۗۗۗۗۗۗۗۗۗۗۗ  ` `L`o`c`k` ` `  pIpnpsp w  wDpeplp w  ` ` `                                                                                                                                                                                  This is the SPACEBAR...                                                         It sort-of reminds us of the space between most users ears.                                                                                                     (Attempts at Humor may not be appreciated during Learning Curves)                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   