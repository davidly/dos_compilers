� �  �                                                                                 ������������������������������������������������������������������������������  �             ����������������������������������������������������           �  �             � Bored of the Look and Feel Police ?              �           �  �             � Or Tired of Eating Your Own Cooking ?            �           �  �             � Log On Today & Check Out What's On The Menu !!!!!�           �  �             ����������������������������������������������������           �  ���������������������������                                                  �  �� Not On The Menu        �          /\              /\              /\      �  ��                        �         /��\            /��\            /��\     �  �� 1. Creamed Silicon     �        /����\          /����\          /����\    �  ��    Chips on Toast      �       /������\        /������\        /������\   �  ��                        �      /Cobalt's\      /��������\      /��������\  �  �� 2. Scrambled           �     /��BOARD���\    /��Bored���\    /��Snorred�\ �  ��    Diskettes           �    /������������\  /������������\  /������������\�  ��                        �    ��������������  ��������������  ���������������  �� 3. Fried Circuits      �    �   �   �   �  �   �    �   �  �   �    �   ��  ��                        �    �  � ?-|�  �  �   �    �   �  �   �    �   ��  �� Exact CRC's Only.      �    ����� ?\ �����  �����    �����  �����    ������  �� We Cannot Make Change. �                                                  �  ���������������������������    COBALT'S HAVEN                                �  ������������������������������������������������������������������������������                                                                                                                                                                                                                                                                                                                                                                                                                 