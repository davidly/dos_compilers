� �  �                                                                                                    -Research Funds are Desperately Needed to Find a Cure                            For Programmer's Insomnia.                                       /\            -Even if I could afford not to I would probably still            //\\            rather do programming all night than Catch Zees.               ///\\\           I would, however, appreciate the opportunity to prove         ////\\\\          or disprove this theory. If you wish to participate in       /////\\\\\         this worthwhile Scientific Experiment and You feel that     ///CANADA\\\        You have received some value from my creations, Please     /������������\       Feel Free To Contribute Whatever Your Conscience Will          �� �� �          Allow. (Preferably money, but anything of value accepted.)     �� �� �                                                                      / / / /b/b/u/c/k/e/l/s/@/m/t/s/./n/e/t/ / / / / / / / / / /B/i/l/l/ /B/u/c/k/e/l/s/,/ /S/t/a/r/v/i/n/g/ /P/r/o/g/r/a/m/m/e/r/ / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / /c///o/ /1/4/ /B/e/r/r/y/d/a/l/e/ /A/v/e/./ / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / /W/i/n/n/i/p/e/g/,/ /M/B/ /R/2/M/1/L/9/ / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / /H/e/r/e/ /I/ / / / / / / / / / / / / / / / / / / / / / / /$/$/$/$/$/$/$/$/$/$/ / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / /�/�/�/�/�/�/�/�/�/�/ / / / / / / / / / / / / / / / / / / /�/�/�/�/�/�/�/�/�/�/ / / / /�/�/�/�/�/ / / / / /�/�/�/ / / / / / / / / / / / / / / / / / / / / / / / /�/�/�/�/�/�/�/�/�/�/ / / / / / / / / / / / / / / / / / / /�/�/�/�/�/�/�/�/�/�/ / / / /�/ / / /�/ / / / / / /�/ / / / / / / / / / /M/a/n/i/t/o/b/a/ / /_/_/_/_/_/�/�/�/�/�/�/�/�/�/�/_/_/_/_/_/C/o/m/e/ / / / / / /_/_/_/_/�/�/�/�/�/�/�/�/�/�/_/_/_/_/�/�/�/�/�/�/�/�/�/�/�/�/�/ / / / / / / / / /�/�/�/�/�/�/�/�/�/�/ / / / / /�/�/�/�/�/�/�/�/�/�/ / / / / /�/�/�/�/�/�/�/�/�/�/ / / / /�/�/�/�/�/�/�/�/�/�/ / / / /�/�/�/�/�/�/�/�/�/�/�/�/�/ / / / / / / / / / / /O/ / / / /O/ / / / / / / / / /O/ / / / /O/ / / / / / / / / /O/ / / / /O/ / / / / / / / /O/ / / / /O/ / / / / / / / / /O/ / / / /O/ / / / /�/ / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / / /N/o/t/e/:/ /I/t/ /i/s/ /o/k/ /t/o/ /m/a/i/l/ /c/a/s/h/,/ /b/u/t/ /d/o/ /n/o/t/ /s/e/n/d/ /c/a/r/s/ /o/r/ /l/i/v/e/s/t/o/c/k/ /t/h/r/o/u/g/h/ /t/h/e/ /m/a/i/l/./� �  �